library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library work;
use work.configuration_pack.all;

entity top_assembler_tb is
--  Port ( );
end top_assembler_tb;

architecture Behavioral of top_assembler_tb is
    component rounding_bits_generator is
      Port ( 
        clk: in std_logic;
        random_rounding_bits: out rounding_bits;
        done: out std_logic
      );
    end component;
    
    
    component MMSU_1 is
      Port ( 
        weight_matrix : in layer_1_w;
        input_vector : in layer_1_in;
        bias_vector: in layer_1_b;
        reset: in std_logic;
        clk: in std_logic;
        random_rounding_bits: in rounding_bits;
        done: out std_logic;
        result : out layer_1_out
      );
    end component;
    
    component VRELU_2 is
      Port ( 
        input: in layer_2_in;
        reset: in std_logic;
        clk: in std_logic;
        done: out std_logic;
        result: out layer_2_out
      );
    end component;
    
    component MMSU_3 is
      Port ( 
        weight_matrix : in layer_3_w;
        input_vector : in layer_3_in;
        bias_vector: in layer_3_b;
        reset: in std_logic;
        clk: in std_logic;
        random_rounding_bits: in rounding_bits;
        done: out std_logic;
        result : out layer_3_out
      );
    end component;
    
    component VRELU_4 is
      Port ( 
        input: in layer_4_in;
        reset: in std_logic;
        clk: in std_logic;
        done: out std_logic;
        result: out layer_4_out
      );
    end component;
    
    component MMSU_5 is
      Port ( 
        weight_matrix : in layer_5_w;
        input_vector : in layer_5_in;
        bias_vector: in layer_5_b;
        reset: in std_logic;
        clk: in std_logic;
        random_rounding_bits: in rounding_bits;
        done: out std_logic;
        result : out layer_5_out
      );
    end component;
    
    component VRELU_6 is
      Port ( 
        input: in layer_6_in;
        reset: in std_logic;
        clk: in std_logic;
        done: out std_logic;
        result: out layer_6_out
      );
    end component;
        
    signal random_rounding_bits: rounding_bits;
    signal clk: std_logic := '0';
    signal generator_done: std_logic;
    signal layer_0_output: layer_0_out;
    
    signal mmsu_1_weight_matrix: layer_1_w;
    signal mmsu_1_bias_vector: layer_1_b;
    signal layer_1_reset: std_logic := '0';
    signal layer_1_done: std_logic := '0';
    signal layer_1_output: layer_1_out; 
    
    signal layer_2_output: layer_2_out;
    signal layer_2_reset, layer_2_done: std_logic;
    
    signal mmsu_3_weight_matrix: layer_3_w;
    signal mmsu_3_bias_vector: layer_3_b;
    signal layer_3_reset: std_logic := '0';
    signal layer_3_done: std_logic := '0';
    signal layer_3_output: layer_3_out;
    
    signal layer_4_output: layer_4_out;
    signal layer_4_reset, layer_4_done: std_logic;
    
    signal mmsu_5_weight_matrix: layer_5_w;
    signal mmsu_5_bias_vector: layer_5_b;
    signal layer_5_reset: std_logic := '0';
    signal layer_5_done: std_logic := '0';
    signal layer_5_output: layer_5_out;
    
    signal layer_6_output: layer_6_out;
    signal layer_6_reset, layer_6_done: std_logic;
    
begin

    layer_2_reset <= not(layer_1_done);
    layer_3_reset <= not(layer_2_done);
    layer_4_reset <= not(layer_3_done);
    layer_5_reset <= not(layer_4_done);
    layer_6_reset <= not(layer_5_done);
    
    GENERATOR: rounding_bits_generator port map(clk => clk, random_rounding_bits => random_rounding_bits, done => generator_done);

    TEST_MMSU_1: MMSU_1 port map(weight_matrix => mmsu_1_weight_matrix, input_vector => layer_0_output, 
                         bias_vector => mmsu_1_bias_vector, reset => layer_1_reset, clk => clk, 
                         random_rounding_bits => random_rounding_bits, done => layer_1_done, 
                         result => layer_1_output);
                         
    TEST_VRELU_2: VRELU_2 port map(input => layer_1_output, reset => layer_2_reset, clk => clk, 
                                     done => layer_2_done, result => layer_2_output);
                                     
    TEST_MMSU_3: MMSU_3 port map(weight_matrix => mmsu_3_weight_matrix, input_vector => layer_2_output, 
                         bias_vector => mmsu_3_bias_vector, reset => layer_3_reset, clk => clk, 
                         random_rounding_bits => random_rounding_bits, done => layer_3_done, 
                         result => layer_3_output);
                         
    TEST_VRELU_4: VRELU_4 port map(input => layer_3_output, reset => layer_4_reset, clk => clk, 
                                     done => layer_4_done, result => layer_4_output);
                                     
    TEST_MMSU_5: MMSU_5 port map(weight_matrix => mmsu_5_weight_matrix, input_vector => layer_4_output, 
                         bias_vector => mmsu_5_bias_vector, reset => layer_5_reset, clk => clk, 
                         random_rounding_bits => random_rounding_bits, done => layer_5_done, 
                         result => layer_5_output);
                         
    TEST_VRELU_6: VRELU_6 port map(input => layer_5_output, reset => layer_6_reset, clk => clk, 
                                     done => layer_6_done, result => layer_6_output);
                         
                         
            
            
    layer_0_output <= ("0000100010101011","1111111001000111","1111101010111110");
                                     
    
    mmsu_1_weight_matrix <= (("0000000001100000","1111111011000011","0000000001010111"),
("0000000010010111","1111111100010000","0000000010000001"),
("0000000000011100","1111111100111010","1111111100111101"),
("1111111100000100","0000000001100100","0000000010110000"),
("1111111011010101","0000000001011110","0000000000101010"),
("0000000011001111","1111111010101001","0000000000000111"),
("1111110111111011","1111111011001010","1111111100101100"),
("0000000000101100","1111111001010101","0000000010111111"),
("0000000011001110","0000000011000111","1111111110010001"),
("1111110101111010","0000000001001010","1111111011100101"),
("0000000100001111","1111111100100111","1111111001101111"),
("1111111101010000","0000000001111101","0000000000010101"),
("0000000100111010","0000000001111101","1111111111001100"),
("1111111110110001","1111111001111001","1111111111101101"),
("1111111000111101","1111111111010110","0000000010011001"),
("1111111111100000","0000000001000010","1111111111100011"));
    
    
    mmsu_1_bias_vector <=  ("0000000011001000","1111111101001011","1111111100100100",
"1111111110011111","0000000110000010","1111111100100100",
"0000000001011011","1111111111111111","0000000101100010",
"0000000111101011","0000000010110111","0000000011110100",
"1111111111101111","1111111100101100","1111110110010100",
"0000000000100001");


    mmsu_3_weight_matrix <= (("1111111111111010","1111111100110110","0000000111011101",
"1111111110100111","0000000100001101","0000000001011011",
"0000000010110001","0000000000100100","0000000010100011",
"0000000100111010","0000000000000000","1111111110111101",
"0000000111000101","1111111100110011","1111111100011110",
"1111111101010111"),
("1111111110010000","0000000110010000","0000000101000010",
"1111111110000101","1111111011100011","0000000101111000",
"1111111111111101","1111111011000000","0000000011001110",
"0000000111000110","1111111110111010","1111111101001000",
"1111111101011101","0000000000100101","1111111100000010",
"1111111101110110"),
("0000000010001010","1111111111101101","1111111111011111",
"0000000001010010","1111111110110100","1111111110110101",
"0000000110000010","1111111001111111","1111111110101101",
"1111111101110011","0000000011110101","0000000010000011",
"0000000011000111","0000000011110100","0000000001011001",
"1111111101100111"),
("1111111001011101","1111111100101101","1111111100010001",
"0000000000001001","1111111111011101","1111111000111001",
"0000000011110011","1111111011001101","0000000011101001",
"1111111110111011","1111111101101000","0000000011011000",
"1111111111001011","0000000010010011","0000000000011001",
"0000000000000001"),
("1111111111111110","1111111100011101","1111111010011100",
"1111111010100010","1111111101001011","1111111101011110",
"0000000110010110","0000000011000101","0000000010011100",
"0000000101000010","1111111011011100","0000000110011001",
"1111111111110011","0000000001100101","1111111001110000",
"1111111011101000"),
("1111111101110010","1111110110111100","0000000000110011",
"0000001000011110","1111111001111111","1111111110100110",
"1111111110001101","0000000110001001","0000000110010011",
"0000000110001101","1111111111010000","0000000001111101",
"1111111101110111","0000000101100001","1111111010110110",
"0000000001110000"),
("0000000010001011","0000000001110111","1111111001010000",
"1111111010101101","1111111101001110","1111111001000101",
"1111111011111110","0000000001010010","0000000001010101",
"1111111110001001","1111111111111001","0000000001111111",
"1111111111110110","1111111010000111","1111111101010101",
"0000000001011011"),
("0000000001110010","1111111000110100","0000000000111110",
"1111111111110110","1111111110100101","0000001010010111",
"0000000111100101","1111111110000000","0000000010101111",
"1111111110000010","1111111110111101","1111111100111111",
"0000000101111101","1111111101001110","1111111001100010",
"1111111111110101"),
("0000000011111110","0000000000100111","0000000001101001",
"0000000011100111","0000000101010110","1111111100100111",
"1111111011011111","0000000000100110","0000000001001011",
"0000000001010011","0000000011011110","0000000011111010",
"0000000000010011","0000000010011100","1111111101111111",
"1111111101011011"),
("0000001010010111","0000000011100111","0000000010101011",
"0000000100110100","0000000011100110","1111111010101001",
"0000000001101001","0000000110000001","0000000100000000",
"0000001000100000","0000000010010000","0000000101110100",
"0000000000110101","0000000111110010","1111111100010101",
"1111111011110101"),
("0000000011100111","1111111100001000","0000000010110100",
"0000000110000110","1111111111100110","0000000011110111",
"0000000110101110","0000000001001100","1111111011110110",
"0000000100101101","0000000000101010","0000000101101000",
"0000000001001000","1111111001110110","0000000000111101",
"1111111111110110"),
("0000000010100101","1111111010111001","0000000011110101",
"0000000000111010","0000000010110110","1111111011101101",
"1111111011111011","0000000011000101","0000000011010101",
"1111111001000001","1111111101100001","0000000000110000",
"1111111110100011","0000000011001101","0000000110101001",
"1111110111111101"),
("1111111110100010","0000000001110101","0000001000101001",
"1111111101000000","1111111011011011","1111111010110010",
"0000000001101010","0000000001001101","0000000001000101",
"0000000001101100","1111111111010101","0000000010000110",
"1111111111010101","0000000110001101","0000000100011100",
"1111111110111101"),
("1111111111010100","0000000001111100","0000000010001101",
"1111111110011001","1111111111011100","0000000010111011",
"1111111110001000","1111111011101011","0000000100100110",
"1111111111110111","0000000000100011","0000000011110100",
"0000000010110110","1111111000001111","0000000001000110",
"1111111101101111"),
("1111111110011110","1111111111010110","0000000010100110",
"1111111101010100","0000000001001001","0000000110010110",
"0000000101010100","0000000011100001","1111111100111111",
"1111111011101011","1111111011010110","0000000011010110",
"0000000010000110","1111111100001011","0000000100100000",
"1111111101100010"),
("0000000011011010","1111110110100010","1111111100111010",
"0000000001101100","0000000000100100","1111111101001110",
"1111111100001101","1111111011111100","1111111101110110",
"1111111001001000","0000001001100111","0000000000001111",
"1111111111010111","1111111100001110","0000000011111001",
"1111111100101101"));


    mmsu_3_bias_vector <= ("0000000100110111","1111111111100111","1111111101000100",
"1111111101110001","0000000011011111","1111111011111111",
"1111111000100100","0000000101101000","0000000000010110",
"1111111110001111","1111111111011011","1111111111001001",
"0000000000101110","1111111111101110","0000000010001111",
"0000000101111010");

    mmsu_5_weight_matrix <= (("1111111101010101","0000000001111101","1111111111100011",
"0000000010110110","0000000010010100","1111111111001101",
"1111111100001011","1111111110011100","0000000101111101",
"0000000011110010","0000000011110010","1111111110101010",
"1111111011110110","1111111011101111","1111111110111011",
"1111111111101100"),
("0000000101111000","0000000101110001","1111111000011111",
"1111111101100011","0000000000011110","1111111101010110",
"1111111101001110","1111111110110000","1111111111111001",
"0000000001111010","1111111001010011","0000000001011101",
"1111111111000001","1111111110111110","1111110110111011",
"1111111101001011"),
("0000000000001011","0000000101110111","0000000100101101",
"1111111101000011","0000001001101111","0000000000001000",
"0000000001001001","0000000011100000","0000000001001000",
"1111111110010101","1111111110010111","1111111000011111",
"1111111111011110","1111111110101110","1111111101111110",
"0000000000001011"));

    mmsu_5_bias_vector <= ("0000000101001101","0000000001001101","0000000010100110");
    
                         
    process
    begin
        clk <= '1';
        wait for 5 ns;
        clk <= '0';
        wait for 5 ns;
    end process;
    
    process
    begin
        layer_1_reset <= '1';
        wait for 10ns;
        layer_1_reset <= '0';
        wait for 1300ns;
    
    end process;
    

end Behavioral;